`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:43:39 12/28/2017 
// Design Name: 
// Module Name:    TC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`define IDLE 2'b00 //
`define LOAD 2'b01
`define CNT  2'b10 // counter
`define INT  2'b11 // interrupt

`define ctrl   mem[0] //���ƼĴ���
`define preset mem[1] //��ֵ�Ĵ���
`define count  mem[2] //����ֵ�Ĵ���

module TC(
    input wire clk,
    input wire reset,
    input wire [31:2] Addr,
    input wire WE, // write enable
    input wire [31:0] Din,
    output wire [31:0] Dout,
    output wire IRQ //interrupt request
    );

	reg [1:0] state;
	reg [31:0] mem [2:0]; // 12B
	
	reg _IRQ;
	assign IRQ = `ctrl[3] & _IRQ;
	
	assign Dout = mem[Addr[3:2]];
	
	wire [31:0] load = Addr[3:2] == 0 ? {28'h0, Din[3:0]} : Din;
	
	integer i;
	always @(posedge clk) begin
		if(reset) begin
			state <= 0; 
			for(i = 0; i < 3; i = i+1) mem[i] <= 0;
			_IRQ <= 0;
		end
		else if(WE) begin
			// $display("%d@: *%h <= %h", $time, {Addr, 2'b00}, load);
			mem[Addr[3:2]] <= load;
		end
		else begin
			case(state)
				`IDLE : if(`ctrl[0]) 
				begin
					state <= `LOAD;
					_IRQ <= 1'b0;
				end
				`LOAD : 
				begin
					`count <= `preset;
					state <= `CNT;
				end
				`CNT  : 
					if(`ctrl[0]) 
					begin
						if(`count > 1) 
							`count <= `count-1;
						else begin
							`count <= 0;
							state <= `INT;
							_IRQ <= 1'b1;
						end
					end
					else 
						state <= `IDLE;
				default : begin
					if(`ctrl[2:1] == 2'b00) 
						`ctrl[0] <= 1'b0;
					else 
						_IRQ <= 1'b0;
					state <= `IDLE;//һ��ִ��
				end
			endcase
		end
	end

endmodule
